`timescale 1ns / 1ps

module tb_TOP_AILayerNorm ();
	reg						i_clk;
	reg						i_rstn;
	reg						i_start;
//	reg	 		[4095:0] 	i_x;
	reg	 		[191:0] 	i_x;
	reg		  	[  7:0] 	i_inv_n;
	reg  		[  1:0] 	i_alpha;
//	reg  		[  7:0] 	i_beta;
//	reg	 		[  7:0]		i_gamma;

	reg  signed	[ 191:0] 	i_beta;
	reg	 signed	[ 191:0]	i_gamma;

//	reg  signed	[4095:0] 	i_beta;
//	reg	 signed	[4095:0]	i_gamma;

	
	wire 					o_done;
	wire signed	[  7:0]		o_AILayerNorm;

	
	always #5 i_clk = ~i_clk;



	TOP_AILayerNorm #(
		.DATA_WIDTH (192)
	)
	u_TOP_AILayerNorm (
		.i_clk(i_clk),
		.i_rstn(i_rstn),
		.i_start(i_start),
		.i_x(i_x),
		.i_inv_n(i_inv_n),
		.i_alpha(i_alpha),
		.i_beta(i_beta),
		.i_gamma(i_gamma),
		.o_done(o_done),
		.o_AILayerNorm(o_AILayerNorm)
	);


	initial 
	begin
		i_clk = 1'd0;		i_rstn = 1'd0;		i_start =  1'd0;	i_x = 192'd0;	
		i_inv_n = 8'd0;		i_alpha = 2'd0;	// 	i_gamma = 8'd0;		i_beta = 8'd0;	
												i_gamma = 192'sd0;	i_beta = 192'sd0;
										//		i_gamma = 4096'sd0;	i_beta = 4096'sd0;
			

		#1 i_rstn = 1'd1;	 #1 i_rstn = 1'd0;	 #4 i_rstn = 1'd1;

		#4 i_start = 1'd1;		i_alpha = 2'd2;		i_inv_n = 8'd32;	//i_gamma = 8'd100;		i_beta = 8'd10;


//  		   i_x = 192'hAC_2F_75_C0_43_FB_C3_67_09_D3_15_F2_24_57_46_D8_58_8C_3A_C1_E6_27_57_AE;

  		   // 192'd172_47_117_192_67_251_195_103_9_211_21_242_36_87_70_216_88_140_58_193_230_39_87_174

//  		   i_x = 320'h00_00_00_00_00_00_00_00_82_82_82_82_82_82_82_82_21_C5_E8_F9_49_B6_1A_F8_00_FF_00_FF_00_FF_00_FF_00_24_48_6C_90_B4_D8_FC;

  		   // 320'd0_0_0_0_0_0_0_0_130_130_130_130_130_130_130_130_33_197_232_249_73_182_26_248_0_255_0_255_0_255_0_255_0_36_72_108_144_180_216_252;


//			i_x = 1024'hAC_2F_75_C0_43_FB_C3_67_09_D3_15_F2_24_57_46_D8_58_8C_3A_C1_E6_27_57_AE_58_51_A5_19_4D_48_09_94_73_D0_F3_C5_FE_4F_AF_C0_52_63_D8_B1_F3_1D_93_93_8E_A7_20_C1_09_B9_7F_20_1F_CA_F4_97_A3_FE_CB_72_B7_1C_22_80_80_A4_35_85_26_E8_F4_11_4F_84_69_2A_BA_1F_78_01_41_E7_A9_39_23_66_77_0B_AE_52_5B_80_8E_63_35_8C_79_AA_54_CB_44_06_C4_2F_7F_F4_83_CC_64_B4_E8_4E_8F_94_E3_BA_17_CF_8D_75_55_30_31_45;
// 1024'd172_47_117_192_67_251_195_103_9_211_21_242_36_87_70_216_88_140_58_193_230_39_87_174_88_81_165_25_77_72_9_148_115_208_243_197_254_79_175_192_82_99_216_177_243_29_147_147_142_167_32_193_9_185_127_32_31_202_244_151_163_254_203_114_183_28_34_128_128_164_53_133_38_232_244_17_79_132_105_42_186_31_120_1_65_231_169_57_35_102_119_11_174_82_91_128_142_99_53_140_121_170_84_203_68_6_196_47_127_244_131_204_100_180_232_78_143_148_227_186_23_207_141_117_85_48_49_69

	//	i_x = 4096'h7C_63_8B_3D_8F_79_51_8F_3E_8C_86_8F_A5_52_29_8D_4A_66_7F_69_62_6C_95_CD_66_51_A4_78_A4_74_6D_AB_92_C6_77_7F_7D_82_EF_5A_A4_97_8D_7C_B0_AA_6A_82_8A_B4_B0_92_79_7F_BD_78_92_62_8C_21_62_6C_79_6A_50_D9_5E_8F_9E_6F_AD_2B_82_7B_73_C1_B4_8A_B0_5F_9B_95_36_66_8A_2E_AE_70_9A_74_A8_AE_65_EE_7A_BB_58_7A_50_5E_66_65_B2_B2_77_6B_46_68_79_53_63_7F_47_4F_AB_6C_B1_AD_8D_79_D6_37_6B_14_8D_5A_9B_C5_A1_87_61_BE_AF_E9_84_78_7F_64_85_88_D9_34_61_66_65_68_99_7A_51_AF_50_98_79_84_5F_34_5C_4A_29_A1_79_7E_93_77_CB_9A_46_01_A7_41_6B_73_82_43_70_65_83_9C_BE_70_8F_89_92_9F_16_37_BC_59_B6_D2_8F_AB_66_35_61_8A_7D_54_5E_8E_80_CD_BA_94_38_7B_D4_43_65_46_7F_56_81_31_8C_50_7C_F4_88_A5_B3_48_54_7D_7D_75_7F_D8_7E_9F_53_1A_59_6A_82_C4_A1_8E_7B_53_55_97_83_63_90_6C_63_24_E2_B0_55_8D_8A_93_54_82_6A_85_81_81_81_45_A3_A7_27_82_A4_4A_52_6B_2E_96_88_8C_62_67_80_84_7C_6C_91_64_A4_89_38_A6_62_BC_75_64_30_7D_38_6A_6C_2A_B3_78_7B_9A_3E_82_5D_51_8A_83_14_84_B2_6D_36_6F_64_67_80_82_99_8F_A0_B6_49_5E_78_93_8A_B8_AE_87_A5_AF_1F_58_94_C4_9B_37_96_67_9F_B3_9F_5F_39_7E_78_94_75_A3_91_61_6D_61_84_A7_C0_31_48_7D_59_A6_7E_51_A2_64_39_4C_7F_9C_9C_7A_8F_4F_C7_A6_C7_9E_C6_76_AE_93_8F_A0_82_92_B6_5A_28_5F_B4_77_81_26_C6_A2_64_4E_37_7F_93_A7_B4_0A_BC_A1_8D_A1_48_A9_37_78_9E_56_78_BA_11_5E_CE_82_BF_75_90_C7_36_59_C7_64_BA_72_60_6B_62_5F_56_92_9C_6C_7A_5E_B9_5E_A0_7C_83_6B_30_85_94_9B_6C_5A_57_AE_8E_BD_A6_82_82_6C_CE_89_6E_4B_71_BE_58_61_9C_30_5B_83_7E_C2_51_9A_9F_BB_84_62_92_9E_98_62_81_A7_62_62_A4_75_33_57_AB_6E_31_2F_8F_98_9A_D4_65_8A_72_82_5B_57_6D_49_7F_9A_6B_2B_9B_A4;


	i_x = 192'h7C_63_8B_3D_8F_79_51_8F_3E_8C_86_8F_A5_52_29_8D_4A_66_7F_69_62_6C_95_CD;
	


	//	i_gamma = 4096'h70_57_58_6C_58_57_55_53_5B_56_59_5B_52_52_5E_58_5A_56_5D_53_5D_58_59_5C_49_59_68_58_4F_5E_58_5A_4E_5A_5D_58_5B_5A_67_5F_65_57_51_55_5B_5D_56_5C_5C_56_4B_57_57_5B_6C_5C_56_56_5C_60_57_5A_5A_60_58_52_51_54_60_57_55_53_59_52_58_56_56_68_5D_5B_56_55_51_55_5D_58_53_58_53_50_5D_5B_5F_57_56_57_5F_5B_59_50_58_5A_57_56_56_59_60_58_52_57_52_5B_56_56_5D_59_5E_5C_59_59_5E_68_54_5A_5D_5A_4F_58_5E_55_4F_62_6B_61_57_5B_58_59_5B_58_5A_59_69_55_59_58_67_54_5D_5B_50_53_5E_59_5D_55_5D_5C_56_60_59_5E_5A_53_5B_54_62_58_58_5E_4E_50_5F_51_5C_59_57_5E_55_5D_59_5B_5A_5A_54_59_59_52_4F_5A_55_58_58_5B_57_5D_5F_52_5D_55_52_54_5E_5F_5B_5B_52_4F_59_57_5A_57_5C_59_65_5A_56_5B_54_5E_59_59_5E_5C_56_56_57_56_59_5E_68_05_5E_5C_5A_4F_5A_64_59_58_5A_59_53_53_5B_50_57_5E_57_5C_52_4D_57_5B_5D_6E_51_5D_54_54_5E_58_54_56_5D_5E_4F_58_51_58_65_58_5E_52_52_5C_58_57_53_60_5C_54_00_59_5B_59_61_5C_5B_4B_55_64_55_4E_5B_59_5F_57_58_61_57_5E_61_4B_51_61_62_58_54_56_5C_58_4D_52_5E_5E_53_5A_5B_53_68_5E_66_57_66_4B_5C_5D_5A_54_56_57_66_56_7D_58_59_50_5A_55_5B_5A_5B_5A_57_5C_5B_57_5E_72_65_5B_5A_55_56_55_53_56_59_59_5A_56_5B_53_55_59_63_5C_5A_51_61_65_56_39_5D_5B_59_57_53_5F_56_58_58_5C_54_58_5A_54_56_51_5B_54_5D_58_5B_59_52_6E_58_59_60_66_59_55_60_56_54_5F_7F_4E_58_57_55_57_5C_5F_61_53_5D_56_00_59_5C_53_55_55_54_66_5A_59_5A_5A_5A_6B_52_52_58_6B_4B_53_55_5E_59_5A_57_53_42_58_62_55_5F_5E_74_57_58_5D_52_60_57_53_55_5B_58_5C_51_56_48_58_54_60_5A_5E_57_54_5A_5A_58_53_5B_55_5C_5B_58_59_58_77_75_60_5D_5E_59_55_60_54_54_78_5B_70_52_51_52_59_5E_52_5A_57_4F_3F_58_53_54_59;

	i_gamma = 192'h70_57_58_6C_58_57_55_53_5B_56_59_5B_52_52_5E_58_5A_56_5D_53_5D_58_59_5C;


	//	i_beta = 4096'h68_08_00_0E_07_E9_1D_E5_F0_03_E4_36_DF_D9_12_D7_DC_F5_12_D4_FC_DF_0E_F2_BA_F6_FC_DD_3A_FB_28_FD_D1_D9_0B_F3_F9_F2_08_B1_19_07_D6_04_E1_F7_13_EA_E9_08_34_D6_10_0E_E8_EE_E4_E4_11_14_E7_F5_07_F9_F5_D2_DF_F7_F9_E0_10_D3_F1_DA_D9_F7_0D_CF_01_C4_D7_DF_02_C6_02_FE_31_DF_E4_E2_15_08_EE_EC_16_13_E7_E8_0F_1D_FB_E2_F2_12_05_06_07_05_18_ED_1F_07_04_2F_2F_01_1B_0F_0C_E8_EC_12_28_16_F4_13_F6_F0_E6_FB_D7_0A_02_D0_1A_16_0A_E8_D9_E5_10_06_05_2E_ED_F3_DE_DC_11_1C_FC_03_1C_E4_04_F5_09_08_E8_EE_E9_2B_FB_27_EF_06_03_EC_14_0D_31_22_1E_31_01_1C_12_05_EC_F6_E7_FC_DD_F5_F5_03_F6_16_D3_E2_0A_19_F8_01_E5_F4_F4_34_13_0D_D9_FB_07_F4_E4_01_24_3C_FD_EF_02_CD_1E_2C_F6_1A_E6_18_17_E8_F3_01_01_F1_CA_D8_00_F7_EE_FC_FE_36_00_18_F8_1F_EB_10_E5_CD_D5_0C_ED_27_E7_E7_E6_F9_1B_05_05_1B_00_F2_04_03_2D_FA_19_E6_FA_F0_C7_01_06_D9_CF_F4_18_0F_E8_13_F9_1B_16_0F_DF_1E_0F_0E_14_EA_03_40_F3_EF_F2_F0_04_D9_CF_13_13_C7_1B_24_2C_09_07_FD_F1_04_0D_B9_1E_0A_FD_0B_2B_0C_E8_FC_C8_25_F7_08_E9_F1_04_0A_FD_0C_CC_FB_10_CA_FA_0E_E6_31_2A_D7_09_FC_F1_13_15_1A_0F_28_DA_F0_FE_F9_E2_F6_F7_DF_13_F8_0D_0F_EE_F8_E5_F8_34_18_F4_05_FE_20_FB_14_F6_05_10_EE_F8_FF_F0_FA_1E_81_02_14_04_E8_EB_0C_F4_14_0E_FA_FE_04_D8_DF_F3_13_E9_E6_36_E3_15_F5_D4_14_15_E7_01_1A_02_24_FE_07_DC_19_E8_EE_E3_17_F3_ED_DE_02_1C_23_E0_13_FB_F0_F8_FD_EA_0B_0C_04_11_D6_F6_13_D2_10_25_22_DF_18_B7_D0_D4_FB_FA_0D_21_25_67_EE_08_DF_0E_E9_16_FF_F0_EA_DB_00_EF_E2_F5_F0_F1_EF_DA_1F_D6_1F_F2_DF_0F_01_11_07_00_F4_01_D4_07_0E_1A_02_EE_FF_21_0B_F6_15_F4_DE_F3_FB_2F_19_FC_02_C4_E5_D0_DE_C8_1A_E5_04_FC_15_36_DE_F6_28_06_0E;

	
	i_beta = 192'h68_08_00_0E_07_E9_1D_E5_F0_03_E4_36_DF_D9_12_D7_DC_F5_12_D4_FC_DF_0E_F2;


		end		   

endmodule
